`define READ_IDLE		2'b00
`define READ_HIT		2'b01
`define READ_STALL		2'b10
`define READ_CHECK		2'b11

module cache_read_sm(
	clk,
	rst,
	rd_en,
	hit,
	mem_done,
	read_state
);

	input clk;
	input rst;
	input rd_en;
	input hit;
	input mem_done;
	output reg [1:0] read_state;

	always @(posedge clk)begin
		if(rst)
			read_state <= `READ_IDLE;
		else
			case(read_state)
				`READ_IDLE: 
					read_state <= rd_en? (hit? `READ_HIT : `READ_STALL) : `READ_IDLE;
				`READ_HIT: 
					read_state <= rd_en? (hit? `READ_HIT : `READ_STALL) : `READ_IDLE;
				`READ_STALL:
					read_state <= (mem_done)? (hit? `READ_HIT : `READ_CHECK) : `READ_STALL;
				`READ_CHECK:
					read_state <= hit? `READ_HIT : `READ_STALL;
				default: 
					read_state <= `READ_IDLE;
			endcase
	end
endmodule
